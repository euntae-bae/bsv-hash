package Tb;

import StmtFSM::*;
import Connectable::*;
import ClientServer::*;

(* synthesize *)
module mkTb(Empty);

endmodule

endpackage