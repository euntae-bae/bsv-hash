package fnlorem;

function Bit#(32) fn_mem_read(Bit#(64) addr);
	return case (addr)
		'h0000000000000000: return 'h4c6f7265;
		'h0000000000000004: return 'h6d206970;
		'h0000000000000008: return 'h73756d20;
		'h000000000000000c: return 'h646f6c6f;
		'h0000000000000010: return 'h72207369;
		'h0000000000000014: return 'h7420616d;
		'h0000000000000018: return 'h65742c20;
		'h000000000000001c: return 'h636f6e73;
		'h0000000000000020: return 'h65637465;
		'h0000000000000024: return 'h74757220;
		'h0000000000000028: return 'h61646970;
		'h000000000000002c: return 'h69736369;
		'h0000000000000030: return 'h6e672065;
		'h0000000000000034: return 'h6c69742e;
		'h0000000000000038: return 'h204d6175;
		'h000000000000003c: return 'h72697320;
		'h0000000000000040: return 'h63757273;
		'h0000000000000044: return 'h75732069;
		'h0000000000000048: return 'h7073756d;
		'h000000000000004c: return 'h20616320;
		'h0000000000000050: return 'h6a757374;
		'h0000000000000054: return 'h6f207665;
		'h0000000000000058: return 'h73746962;
		'h000000000000005c: return 'h756c756d;
		'h0000000000000060: return 'h20646170;
		'h0000000000000064: return 'h69627573;
		'h0000000000000068: return 'h2e20446f;
		'h000000000000006c: return 'h6e656320;
		'h0000000000000070: return 'h73616769;
		'h0000000000000074: return 'h74746973;
		'h0000000000000078: return 'h206d6f6c;
		'h000000000000007c: return 'h6c697320;
		'h0000000000000080: return 'h74656d70;
		'h0000000000000084: return 'h6f722e20;
		'h0000000000000088: return 'h496e7465;
		'h000000000000008c: return 'h67657220;
		'h0000000000000090: return 'h636f6e73;
		'h0000000000000094: return 'h65637465;
		'h0000000000000098: return 'h74757220;
		'h000000000000009c: return 'h69707375;
		'h00000000000000a0: return 'h6d207465;
		'h00000000000000a4: return 'h6c6c7573;
		'h00000000000000a8: return 'h2c207365;
		'h00000000000000ac: return 'h6420636f;
		'h00000000000000b0: return 'h6e76616c;
		'h00000000000000b4: return 'h6c697320;
		'h00000000000000b8: return 'h66656c69;
		'h00000000000000bc: return 'h7320656c;
		'h00000000000000c0: return 'h65696665;
		'h00000000000000c4: return 'h6e642061;
		'h00000000000000c8: return 'h742e2055;
		'h00000000000000cc: return 'h74206575;
		'h00000000000000d0: return 'h206d6920;
		'h00000000000000d4: return 'h656c6974;
		'h00000000000000d8: return 'h2e205375;
		'h00000000000000dc: return 'h7370656e;
		'h00000000000000e0: return 'h64697373;
		'h00000000000000e4: return 'h65206772;
		'h00000000000000e8: return 'h61766964;
		'h00000000000000ec: return 'h61206661;
		'h00000000000000f0: return 'h75636962;
		'h00000000000000f4: return 'h75732074;
		'h00000000000000f8: return 'h656c6c75;
		'h00000000000000fc: return 'h7320636f;
		'h0000000000000100: return 'h6e736563;
		'h0000000000000104: return 'h74657475;
		'h0000000000000108: return 'h72207465;
		'h000000000000010c: return 'h6d707573;
		'h0000000000000110: return 'h2e204165;
		'h0000000000000114: return 'h6e65616e;
		'h0000000000000118: return 'h206e6563;
		'h000000000000011c: return 'h206c6967;
		'h0000000000000120: return 'h756c6120;
		'h0000000000000124: return 'h76656c20;
		'h0000000000000128: return 'h61726375;
		'h000000000000012c: return 'h20756c74;
		'h0000000000000130: return 'h72696369;
		'h0000000000000134: return 'h65732066;
		'h0000000000000138: return 'h61756369;
		'h000000000000013c: return 'h62757320;
		'h0000000000000140: return 'h6e6f6e20;
		'h0000000000000144: return 'h65752070;
		'h0000000000000148: return 'h75727573;
		'h000000000000014c: return 'h2e20496e;
		'h0000000000000150: return 'h74656765;
		'h0000000000000154: return 'h72207465;
		'h0000000000000158: return 'h6d706f72;
		'h000000000000015c: return 'h2074656c;
		'h0000000000000160: return 'h6c757320;
		'h0000000000000164: return 'h73697420;
		'h0000000000000168: return 'h616d6574;
		'h000000000000016c: return 'h2074696e;
		'h0000000000000170: return 'h63696475;
		'h0000000000000174: return 'h6e74206d;
		'h0000000000000178: return 'h6178696d;
		'h000000000000017c: return 'h75732e20;
		'h0000000000000180: return 'h496e2076;
		'h0000000000000184: return 'h65737469;
		'h0000000000000188: return 'h62756c75;
		'h000000000000018c: return 'h6d206e69;
		'h0000000000000190: return 'h6268206d;
		'h0000000000000194: return 'h65747573;
		'h0000000000000198: return 'h2c206163;
		'h000000000000019c: return 'h20706f73;
		'h00000000000001a0: return 'h75657265;
		'h00000000000001a4: return 'h206d6574;
		'h00000000000001a8: return 'h75732062;
		'h00000000000001ac: return 'h6c616e64;
		'h00000000000001b0: return 'h69742076;
		'h00000000000001b4: return 'h69746165;
		'h00000000000001b8: return 'h2e204c6f;
		'h00000000000001bc: return 'h72656d20;
		'h00000000000001c0: return 'h69707375;
		'h00000000000001c4: return 'h6d20646f;
		'h00000000000001c8: return 'h6c6f7220;
		'h00000000000001cc: return 'h73697420;
		'h00000000000001d0: return 'h616d6574;
		'h00000000000001d4: return 'h2c20636f;
		'h00000000000001d8: return 'h6e736563;
		'h00000000000001dc: return 'h74657475;
		'h00000000000001e0: return 'h72206164;
		'h00000000000001e4: return 'h69706973;
		'h00000000000001e8: return 'h63696e67;
		'h00000000000001ec: return 'h20656c69;
		'h00000000000001f0: return 'h742e2049;
		'h00000000000001f4: return 'h6e746567;
		'h00000000000001f8: return 'h65722065;
		'h00000000000001fc: return 'h6c656d65;
		'h0000000000000200: return 'h6e74756d;
		'h0000000000000204: return 'h20657261;
		'h0000000000000208: return 'h74206574;
		'h000000000000020c: return 'h20736f64;
		'h0000000000000210: return 'h616c6573;
		'h0000000000000214: return 'h20736f6c;
		'h0000000000000218: return 'h6c696369;
		'h000000000000021c: return 'h74756469;
		'h0000000000000220: return 'h6e2e204e;
		'h0000000000000224: return 'h756c6c61;
		'h0000000000000228: return 'h6d206567;
		'h000000000000022c: return 'h6574206f;
		'h0000000000000230: return 'h64696f20;
		'h0000000000000234: return 'h6c656374;
		'h0000000000000238: return 'h75732e20;
		'h000000000000023c: return 'h45746961;
		'h0000000000000240: return 'h6d206961;
		'h0000000000000244: return 'h63756c69;
		'h0000000000000248: return 'h73206f72;
		'h000000000000024c: return 'h6369206c;
		'h0000000000000250: return 'h69626572;
		'h0000000000000254: return 'h6f2e2056;
		'h0000000000000258: return 'h6976616d;
		'h000000000000025c: return 'h75732061;
		'h0000000000000260: return 'h6c697175;
		'h0000000000000264: return 'h65742061;
		'h0000000000000268: return 'h6e746520;
		'h000000000000026c: return 'h65742064;
		'h0000000000000270: return 'h75692061;
		'h0000000000000274: return 'h6c697175;
		'h0000000000000278: return 'h65742c20;
		'h000000000000027c: return 'h65752065;
		'h0000000000000280: return 'h6c656d65;
		'h0000000000000284: return 'h6e74756d;
		'h0000000000000288: return 'h206d6173;
		'h000000000000028c: return 'h73612073;
		'h0000000000000290: return 'h6f64616c;
		'h0000000000000294: return 'h65732e20;
		'h0000000000000298: return 'h50656c6c;
		'h000000000000029c: return 'h656e7465;
		'h00000000000002a0: return 'h73717565;
		'h00000000000002a4: return 'h20736f64;
		'h00000000000002a8: return 'h616c6573;
		'h00000000000002ac: return 'h20657374;
		'h00000000000002b0: return 'h2061206e;
		'h00000000000002b4: return 'h69736c20;
		'h00000000000002b8: return 'h636f6e73;
		'h00000000000002bc: return 'h65637465;
		'h00000000000002c0: return 'h7475722c;
		'h00000000000002c4: return 'h20696420;
		'h00000000000002c8: return 'h706f7274;
		'h00000000000002cc: return 'h7469746f;
		'h00000000000002d0: return 'h72206d61;
		'h00000000000002d4: return 'h73736120;
		'h00000000000002d8: return 'h70726574;
		'h00000000000002dc: return 'h69756d2e;
		default: return 0;
	endcase;
endfunction

endpackage