package Jhash;

interface Jhash_IFC;
endinterface

module mkJhash(Jhash_IFC);
endmodule

endpackage