package Tb;

endpackage